LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY nand8 IS
  PORT
  (
    in1  : IN std_logic_vector(7 DOWNTO 0);
    out1 : OUT std_logic_vector(7 DOWNTO 0)
  );
END ENTITY nand8;


architecture genericType of nand8 is
  
begin
  
  
  
end architecture genericType;